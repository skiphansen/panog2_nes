// Based on apu.sv from https://github.com/MiSTer-devel/NES_MiSTer.git

// Copyright (c) 2012-2013 Ludvig Strigeus
// This program is GPL Licensed. See COPYING for the full license.
 

// http://wiki.nesdev.com/w/index.php/APU_Mixer
// I generated three LUT's for each mix channel entry and one lut for the squares, then a
// 282 entry lut for the mix channel. It's more accurate than the original LUT system listed on
// the NesDev page.

module APUMixer (
  input [3:0] square1,
  input [3:0] square2,
  input [3:0] triangle,
  input [3:0] noise,
  input [6:0] dmc,
  output reg [15:0] sample
);


wire [4:0] squares = square1 + square2;
// wire [8:0] mix = tri_lut[triangle] + noise_lut[noise] + dmc_lut[dmc];

reg [5:0] tri_lookup;
reg [3:0] noise_lookup;
reg [6:0] dmc_lookup;
reg [8:0] mix;
reg [15:0] ch1;
reg [15:0] ch2;
reg [16:0] chan_mix;

always @*
  begin
    tri_lookup = 6'd0;

    case (triangle)
        4'd0 : tri_lookup = 6'd0;
        4'd1 : tri_lookup = 6'd3;
        4'd2 : tri_lookup = 6'd7;
        4'd3 : tri_lookup = 6'd11;
        4'd4 : tri_lookup = 6'd15;
        4'd5 : tri_lookup = 6'd19;
        4'd6 : tri_lookup = 6'd23;
        4'd7 : tri_lookup = 6'd27;
        4'd8 : tri_lookup = 6'd31;
        4'd9 : tri_lookup = 6'd35;
        4'd10 : tri_lookup = 6'd39;
        4'd11 : tri_lookup = 6'd43;
        4'd12 : tri_lookup = 6'd47;
        4'd13 : tri_lookup = 6'd51;
        4'd14 : tri_lookup = 6'd55;
        4'd15 : tri_lookup = 6'd59;
    endcase

    case (noise)
        4'd0 : noise_lookup = 6'd0;
        4'd1 : noise_lookup = 6'd2;
        4'd2 : noise_lookup = 6'd5;
        4'd3 : noise_lookup = 6'd8;
        4'd4 : noise_lookup = 6'd10;
        4'd5 : noise_lookup = 6'd13;
        4'd6 : noise_lookup = 6'd16;
        4'd7 : noise_lookup = 6'd18;
        4'd8 : noise_lookup = 6'd21;
        4'd9 : noise_lookup = 6'd24;
        4'd10 : noise_lookup = 6'd26;
        4'd11 : noise_lookup = 6'd29;
        4'd12 : noise_lookup = 6'd32;
        4'd13 : noise_lookup = 6'd34;
        4'd14 : noise_lookup = 6'd37;
        4'd15 : noise_lookup = 6'd40;
    endcase

    case (dmc)
        7'd0 : dmc_lookup = 8'd0;
        7'd1 : dmc_lookup = 8'd1;
        7'd2 : dmc_lookup = 8'd2;
        7'd3 : dmc_lookup = 8'd4;
        7'd4 : dmc_lookup = 8'd5;
        7'd5 : dmc_lookup = 8'd7;
        7'd6 : dmc_lookup = 8'd8;
        7'd7 : dmc_lookup = 8'd10;
        7'd8 : dmc_lookup = 8'd11;
        7'd9 : dmc_lookup = 8'd13;
        7'd10 : dmc_lookup = 8'd14;
        7'd11 : dmc_lookup = 8'd15;
        7'd12 : dmc_lookup = 8'd17;
        7'd13 : dmc_lookup = 8'd18;
        7'd14 : dmc_lookup = 8'd20;
        7'd15 : dmc_lookup = 8'd21;
        7'd16 : dmc_lookup = 8'd23;
        7'd17 : dmc_lookup = 8'd24;
        7'd18 : dmc_lookup = 8'd26;
        7'd19 : dmc_lookup = 8'd27;
        7'd20 : dmc_lookup = 8'd28;
        7'd21 : dmc_lookup = 8'd30;
        7'd22 : dmc_lookup = 8'd31;
        7'd23 : dmc_lookup = 8'd33;
        7'd24 : dmc_lookup = 8'd34;
        7'd25 : dmc_lookup = 8'd36;
        7'd26 : dmc_lookup = 8'd37;
        7'd27 : dmc_lookup = 8'd39;
        7'd28 : dmc_lookup = 8'd40;
        7'd29 : dmc_lookup = 8'd41;
        7'd30 : dmc_lookup = 8'd43;
        7'd31 : dmc_lookup = 8'd44;
        7'd32 : dmc_lookup = 8'd46;
        7'd33 : dmc_lookup = 8'd47;
        7'd34 : dmc_lookup = 8'd49;
        7'd35 : dmc_lookup = 8'd50;
        7'd36 : dmc_lookup = 8'd52;
        7'd37 : dmc_lookup = 8'd53;
        7'd38 : dmc_lookup = 8'd55;
        7'd39 : dmc_lookup = 8'd56;
        7'd40 : dmc_lookup = 8'd57;
        7'd41 : dmc_lookup = 8'd59;
        7'd42 : dmc_lookup = 8'd60;
        7'd43 : dmc_lookup = 8'd62;
        7'd44 : dmc_lookup = 8'd63;
        7'd45 : dmc_lookup = 8'd65;
        7'd46 : dmc_lookup = 8'd66;
        7'd47 : dmc_lookup = 8'd68;
        7'd48 : dmc_lookup = 8'd69;
        7'd49 : dmc_lookup = 8'd70;
        7'd50 : dmc_lookup = 8'd72;
        7'd51 : dmc_lookup = 8'd73;
        7'd52 : dmc_lookup = 8'd75;
        7'd53 : dmc_lookup = 8'd76;
        7'd54 : dmc_lookup = 8'd78;
        7'd55 : dmc_lookup = 8'd79;
        7'd56 : dmc_lookup = 8'd81;
        7'd57 : dmc_lookup = 8'd82;
        7'd58 : dmc_lookup = 8'd83;
        7'd59 : dmc_lookup = 8'd85;
        7'd60 : dmc_lookup = 8'd86;
        7'd61 : dmc_lookup = 8'd88;
        7'd62 : dmc_lookup = 8'd89;
        7'd63 : dmc_lookup = 8'd91;
        7'd64 : dmc_lookup = 8'd92;
        7'd65 : dmc_lookup = 8'd94;
        7'd66 : dmc_lookup = 8'd95;
        7'd67 : dmc_lookup = 8'd96;
        7'd68 : dmc_lookup = 8'd98;
        7'd69 : dmc_lookup = 8'd99;
        7'd70 : dmc_lookup = 8'd101;
        7'd71 : dmc_lookup = 8'd102;
        7'd72 : dmc_lookup = 8'd104;
        7'd73 : dmc_lookup = 8'd105;
        7'd74 : dmc_lookup = 8'd107;
        7'd75 : dmc_lookup = 8'd108;
        7'd76 : dmc_lookup = 8'd110;
        7'd77 : dmc_lookup = 8'd111;
        7'd78 : dmc_lookup = 8'd112;
        7'd79 : dmc_lookup = 8'd114;
        7'd80 : dmc_lookup = 8'd115;
        7'd81 : dmc_lookup = 8'd117;
        7'd82 : dmc_lookup = 8'd118;
        7'd83 : dmc_lookup = 8'd120;
        7'd84 : dmc_lookup = 8'd121;
        7'd85 : dmc_lookup = 8'd123;
        7'd86 : dmc_lookup = 8'd124;
        7'd87 : dmc_lookup = 8'd125;
        7'd88 : dmc_lookup = 8'd127;
        7'd89 : dmc_lookup = 8'd128;
        7'd90 : dmc_lookup = 8'd130;
        7'd91 : dmc_lookup = 8'd131;
        7'd92 : dmc_lookup = 8'd133;
        7'd93 : dmc_lookup = 8'd134;
        7'd94 : dmc_lookup = 8'd136;
        7'd95 : dmc_lookup = 8'd137;
        7'd96 : dmc_lookup = 8'd138;
        7'd97 : dmc_lookup = 8'd140;
        7'd98 : dmc_lookup = 8'd141;
        7'd99 : dmc_lookup = 8'd143;
        7'd100 : dmc_lookup = 8'd144;
        7'd101 : dmc_lookup = 8'd146;
        7'd102 : dmc_lookup = 8'd147;
        7'd103 : dmc_lookup = 8'd149;
        7'd104 : dmc_lookup = 8'd150;
        7'd105 : dmc_lookup = 8'd151;
        7'd106 : dmc_lookup = 8'd153;
        7'd107 : dmc_lookup = 8'd154;
        7'd108 : dmc_lookup = 8'd156;
        7'd109 : dmc_lookup = 8'd157;
        7'd110 : dmc_lookup = 8'd159;
        7'd111 : dmc_lookup = 8'd160;
        7'd112 : dmc_lookup = 8'd162;
        7'd113 : dmc_lookup = 8'd163;
        7'd114 : dmc_lookup = 8'd165;
        7'd115 : dmc_lookup = 8'd166;
        7'd116 : dmc_lookup = 8'd167;
        7'd117 : dmc_lookup = 8'd169;
        7'd118 : dmc_lookup = 8'd170;
        7'd119 : dmc_lookup = 8'd172;
        7'd120 : dmc_lookup = 8'd173;
        7'd121 : dmc_lookup = 8'd175;
        7'd122 : dmc_lookup = 8'd176;
        7'd123 : dmc_lookup = 8'd178;
        7'd124 : dmc_lookup = 8'd179;
        7'd125 : dmc_lookup = 8'd180;
        7'd126 : dmc_lookup = 8'd182;
        7'd127 : dmc_lookup = 8'd183;
    endcase

    mix = tri_lookup + noise_lookup + dmc_lookup;

    // wire [15:0] ch1 = pulse_lut[squares];
    case (squares)
        6'd0 : ch1 = 16'd0;
        6'd1 : ch1 = 16'd763;
        6'd2 : ch1 = 16'd1509;
        6'd3 : ch1 = 16'd2236;
        6'd4 : ch1 = 16'd2947;
        6'd5 : ch1 = 16'd3641;
        6'd6 : ch1 = 16'd4319;
        6'd7 : ch1 = 16'd4982;
        6'd8 : ch1 = 16'd5630;
        6'd9 : ch1 = 16'd6264;
        6'd10 : ch1 = 16'd6883;
        6'd11 : ch1 = 16'd7490;
        6'd12 : ch1 = 16'd8083;
        6'd13 : ch1 = 16'd8664;
        6'd14 : ch1 = 16'd9232;
        6'd15 : ch1 = 16'd9789;
        6'd16 : ch1 = 16'd10334;
        6'd17 : ch1 = 16'd10868;
        6'd18 : ch1 = 16'd11392;
        6'd19 : ch1 = 16'd11905;
        6'd20 : ch1 = 16'd12408;
        6'd21 : ch1 = 16'd12901;
        6'd22 : ch1 = 16'd13384;
        6'd23 : ch1 = 16'd13858;
        6'd24 : ch1 = 16'd14324;
        6'd25 : ch1 = 16'd14780;
        6'd26 : ch1 = 16'd15228;
        6'd27 : ch1 = 16'd15668;
        6'd28 : ch1 = 16'd16099;
        6'd29 : ch1 = 16'd16523;
        6'd30 : ch1 = 16'd16939;
        6'd31 : ch1 = 16'd17348;
    endcase


    // wire [15:0] ch2 = mix_lut[mix];
    case (mix)
        9'd0 : ch2 = 16'd0;
        9'd1 : ch2 = 16'd318;
        9'd2 : ch2 = 16'd635;
        9'd3 : ch2 = 16'd950;
        9'd4 : ch2 = 16'd1262;
        9'd5 : ch2 = 16'd1573;
        9'd6 : ch2 = 16'd1882;
        9'd7 : ch2 = 16'd2190;
        9'd8 : ch2 = 16'd2495;
        9'd9 : ch2 = 16'd2799;
        9'd10 : ch2 = 16'd3101;
        9'd11 : ch2 = 16'd3401;
        9'd12 : ch2 = 16'd3699;
        9'd13 : ch2 = 16'd3995;
        9'd14 : ch2 = 16'd4290;
        9'd15 : ch2 = 16'd4583;
        9'd16 : ch2 = 16'd4875;
        9'd17 : ch2 = 16'd5164;
        9'd18 : ch2 = 16'd5452;
        9'd19 : ch2 = 16'd5739;
        9'd20 : ch2 = 16'd6023;
        9'd21 : ch2 = 16'd6306;
        9'd22 : ch2 = 16'd6588;
        9'd23 : ch2 = 16'd6868;
        9'd24 : ch2 = 16'd7146;
        9'd25 : ch2 = 16'd7423;
        9'd26 : ch2 = 16'd7698;
        9'd27 : ch2 = 16'd7971;
        9'd28 : ch2 = 16'd8243;
        9'd29 : ch2 = 16'd8514;
        9'd30 : ch2 = 16'd8783;
        9'd31 : ch2 = 16'd9050;
        9'd32 : ch2 = 16'd9316;
        9'd33 : ch2 = 16'd9581;
        9'd34 : ch2 = 16'd9844;
        9'd35 : ch2 = 16'd10105;
        9'd36 : ch2 = 16'd10365;
        9'd37 : ch2 = 16'd10624;
        9'd38 : ch2 = 16'd10881;
        9'd39 : ch2 = 16'd11137;
        9'd40 : ch2 = 16'd11392;
        9'd41 : ch2 = 16'd11645;
        9'd42 : ch2 = 16'd11897;
        9'd43 : ch2 = 16'd12147;
        9'd44 : ch2 = 16'd12396;
        9'd45 : ch2 = 16'd12644;
        9'd46 : ch2 = 16'd12890;
        9'd47 : ch2 = 16'd13135;
        9'd48 : ch2 = 16'd13379;
        9'd49 : ch2 = 16'd13622;
        9'd50 : ch2 = 16'd13863;
        9'd51 : ch2 = 16'd14103;
        9'd52 : ch2 = 16'd14341;
        9'd53 : ch2 = 16'd14579;
        9'd54 : ch2 = 16'd14815;
        9'd55 : ch2 = 16'd15050;
        9'd56 : ch2 = 16'd15284;
        9'd57 : ch2 = 16'd15516;
        9'd58 : ch2 = 16'd15747;
        9'd59 : ch2 = 16'd15978;
        9'd60 : ch2 = 16'd16206;
        9'd61 : ch2 = 16'd16434;
        9'd62 : ch2 = 16'd16661;
        9'd63 : ch2 = 16'd16886;
        9'd64 : ch2 = 16'd17110;
        9'd65 : ch2 = 16'd17333;
        9'd66 : ch2 = 16'd17555;
        9'd67 : ch2 = 16'd17776;
        9'd68 : ch2 = 16'd17996;
        9'd69 : ch2 = 16'd18215;
        9'd70 : ch2 = 16'd18432;
        9'd71 : ch2 = 16'd18649;
        9'd72 : ch2 = 16'd18864;
        9'd73 : ch2 = 16'd19078;
        9'd74 : ch2 = 16'd19291;
        9'd75 : ch2 = 16'd19504;
        9'd76 : ch2 = 16'd19715;
        9'd77 : ch2 = 16'd19925;
        9'd78 : ch2 = 16'd20134;
        9'd79 : ch2 = 16'd20342;
        9'd80 : ch2 = 16'd20549;
        9'd81 : ch2 = 16'd20755;
        9'd82 : ch2 = 16'd20960;
        9'd83 : ch2 = 16'd21163;
        9'd84 : ch2 = 16'd21366;
        9'd85 : ch2 = 16'd21568;
        9'd86 : ch2 = 16'd21769;
        9'd87 : ch2 = 16'd21969;
        9'd88 : ch2 = 16'd22169;
        9'd89 : ch2 = 16'd22367;
        9'd90 : ch2 = 16'd22564;
        9'd91 : ch2 = 16'd22760;
        9'd92 : ch2 = 16'd22955;
        9'd93 : ch2 = 16'd23150;
        9'd94 : ch2 = 16'd23343;
        9'd95 : ch2 = 16'd23536;
        9'd96 : ch2 = 16'd23727;
        9'd97 : ch2 = 16'd23918;
        9'd98 : ch2 = 16'd24108;
        9'd99 : ch2 = 16'd24297;
        9'd100 : ch2 = 16'd24485;
        9'd101 : ch2 = 16'd24672;
        9'd102 : ch2 = 16'd24858;
        9'd103 : ch2 = 16'd25044;
        9'd104 : ch2 = 16'd25228;
        9'd105 : ch2 = 16'd25412;
        9'd106 : ch2 = 16'd25595;
        9'd107 : ch2 = 16'd25777;
        9'd108 : ch2 = 16'd25958;
        9'd109 : ch2 = 16'd26138;
        9'd110 : ch2 = 16'd26318;
        9'd111 : ch2 = 16'd26497;
        9'd112 : ch2 = 16'd26674;
        9'd113 : ch2 = 16'd26852;
        9'd114 : ch2 = 16'd27028;
        9'd115 : ch2 = 16'd27203;
        9'd116 : ch2 = 16'd27378;
        9'd117 : ch2 = 16'd27552;
        9'd118 : ch2 = 16'd27725;
        9'd119 : ch2 = 16'd27898;
        9'd120 : ch2 = 16'd28069;
        9'd121 : ch2 = 16'd28240;
        9'd122 : ch2 = 16'd28410;
        9'd123 : ch2 = 16'd28579;
        9'd124 : ch2 = 16'd28748;
        9'd125 : ch2 = 16'd28916;
        9'd126 : ch2 = 16'd29083;
        9'd127 : ch2 = 16'd29249;
        9'd128 : ch2 = 16'd29415;
        9'd129 : ch2 = 16'd29580;
        9'd130 : ch2 = 16'd29744;
        9'd131 : ch2 = 16'd29907;
        9'd132 : ch2 = 16'd30070;
        9'd133 : ch2 = 16'd30232;
        9'd134 : ch2 = 16'd30393;
        9'd135 : ch2 = 16'd30554;
        9'd136 : ch2 = 16'd30714;
        9'd137 : ch2 = 16'd30873;
        9'd138 : ch2 = 16'd31032;
        9'd139 : ch2 = 16'd31190;
        9'd140 : ch2 = 16'd31347;
        9'd141 : ch2 = 16'd31503;
        9'd142 : ch2 = 16'd31659;
        9'd143 : ch2 = 16'd31815;
        9'd144 : ch2 = 16'd31969;
        9'd145 : ch2 = 16'd32123;
        9'd146 : ch2 = 16'd32276;
        9'd147 : ch2 = 16'd32429;
        9'd148 : ch2 = 16'd32581;
        9'd149 : ch2 = 16'd32732;
        9'd150 : ch2 = 16'd32883;
        9'd151 : ch2 = 16'd33033;
        9'd152 : ch2 = 16'd33182;
        9'd153 : ch2 = 16'd33331;
        9'd154 : ch2 = 16'd33479;
        9'd155 : ch2 = 16'd33627;
        9'd156 : ch2 = 16'd33774;
        9'd157 : ch2 = 16'd33920;
        9'd158 : ch2 = 16'd34066;
        9'd159 : ch2 = 16'd34211;
        9'd160 : ch2 = 16'd34356;
        9'd161 : ch2 = 16'd34500;
        9'd162 : ch2 = 16'd34643;
        9'd163 : ch2 = 16'd34786;
        9'd164 : ch2 = 16'd34928;
        9'd165 : ch2 = 16'd35070;
        9'd166 : ch2 = 16'd35211;
        9'd167 : ch2 = 16'd35352;
        9'd168 : ch2 = 16'd35492;
        9'd169 : ch2 = 16'd35631;
        9'd170 : ch2 = 16'd35770;
        9'd171 : ch2 = 16'd35908;
        9'd172 : ch2 = 16'd36046;
        9'd173 : ch2 = 16'd36183;
        9'd174 : ch2 = 16'd36319;
        9'd175 : ch2 = 16'd36456;
        9'd176 : ch2 = 16'd36591;
        9'd177 : ch2 = 16'd36726;
        9'd178 : ch2 = 16'd36860;
        9'd179 : ch2 = 16'd36994;
        9'd180 : ch2 = 16'd37128;
        9'd181 : ch2 = 16'd37261;
        9'd182 : ch2 = 16'd37393;
        9'd183 : ch2 = 16'd37525;
        9'd184 : ch2 = 16'd37656;
        9'd185 : ch2 = 16'd37787;
        9'd186 : ch2 = 16'd37917;
        9'd187 : ch2 = 16'd38047;
        9'd188 : ch2 = 16'd38176;
        9'd189 : ch2 = 16'd38305;
        9'd190 : ch2 = 16'd38433;
        9'd191 : ch2 = 16'd38561;
        9'd192 : ch2 = 16'd38689;
        9'd193 : ch2 = 16'd38815;
        9'd194 : ch2 = 16'd38942;
        9'd195 : ch2 = 16'd39068;
        9'd196 : ch2 = 16'd39193;
        9'd197 : ch2 = 16'd39318;
        9'd198 : ch2 = 16'd39442;
        9'd199 : ch2 = 16'd39566;
        9'd200 : ch2 = 16'd39690;
        9'd201 : ch2 = 16'd39813;
        9'd202 : ch2 = 16'd39935;
        9'd203 : ch2 = 16'd40057;
        9'd204 : ch2 = 16'd40179;
        9'd205 : ch2 = 16'd40300;
        9'd206 : ch2 = 16'd40421;
        9'd207 : ch2 = 16'd40541;
        9'd208 : ch2 = 16'd40661;
        9'd209 : ch2 = 16'd40780;
        9'd210 : ch2 = 16'd40899;
        9'd211 : ch2 = 16'd41017;
        9'd212 : ch2 = 16'd41136;
        9'd213 : ch2 = 16'd41253;
        9'd214 : ch2 = 16'd41370;
        9'd215 : ch2 = 16'd41487;
        9'd216 : ch2 = 16'd41603;
        9'd217 : ch2 = 16'd41719;
        9'd218 : ch2 = 16'd41835;
        9'd219 : ch2 = 16'd41950;
        9'd220 : ch2 = 16'd42064;
        9'd221 : ch2 = 16'd42178;
        9'd222 : ch2 = 16'd42292;
        9'd223 : ch2 = 16'd42406;
        9'd224 : ch2 = 16'd42519;
        9'd225 : ch2 = 16'd42631;
        9'd226 : ch2 = 16'd42743;
        9'd227 : ch2 = 16'd42855;
        9'd228 : ch2 = 16'd42966;
        9'd229 : ch2 = 16'd43077;
        9'd230 : ch2 = 16'd43188;
        9'd231 : ch2 = 16'd43298;
        9'd232 : ch2 = 16'd43408;
        9'd233 : ch2 = 16'd43517;
        9'd234 : ch2 = 16'd43626;
        9'd235 : ch2 = 16'd43735;
        9'd236 : ch2 = 16'd43843;
        9'd237 : ch2 = 16'd43951;
        9'd238 : ch2 = 16'd44058;
        9'd239 : ch2 = 16'd44165;
        9'd240 : ch2 = 16'd44272;
        9'd241 : ch2 = 16'd44378;
        9'd242 : ch2 = 16'd44484;
        9'd243 : ch2 = 16'd44589;
        9'd244 : ch2 = 16'd44695;
        9'd245 : ch2 = 16'd44799;
        9'd246 : ch2 = 16'd44904;
        9'd247 : ch2 = 16'd45008;
        9'd248 : ch2 = 16'd45112;
        9'd249 : ch2 = 16'd45215;
        9'd250 : ch2 = 16'd45318;
        9'd251 : ch2 = 16'd45421;
        9'd252 : ch2 = 16'd45523;
        9'd253 : ch2 = 16'd45625;
        9'd254 : ch2 = 16'd45726;
        9'd255 : ch2 = 16'd45828;
        9'd256 : ch2 = 16'd45929;
        9'd257 : ch2 = 16'd46029;
        9'd258 : ch2 = 16'd46129;
        9'd259 : ch2 = 16'd46229;
        9'd260 : ch2 = 16'd46329;
        9'd261 : ch2 = 16'd46428;
        9'd262 : ch2 = 16'd46527;
        9'd263 : ch2 = 16'd46625;
        9'd264 : ch2 = 16'd46723;
        9'd265 : ch2 = 16'd46821;
        9'd266 : ch2 = 16'd46919;
        9'd267 : ch2 = 16'd47016;
        9'd268 : ch2 = 16'd47113;
        9'd269 : ch2 = 16'd47209;
        9'd270 : ch2 = 16'd47306;
        9'd271 : ch2 = 16'd47402;
        9'd272 : ch2 = 16'd47497;
        9'd273 : ch2 = 16'd47592;
        9'd274 : ch2 = 16'd47687;
        9'd275 : ch2 = 16'd47782;
        9'd276 : ch2 = 16'd47876;
        9'd277 : ch2 = 16'd47970;
        9'd278 : ch2 = 16'd48064;
        9'd279 : ch2 = 16'd48157;
        9'd280 : ch2 = 16'd48250;
        9'd281 : ch2 = 16'd48343;
        9'd282 : ch2 = 16'd48436;
        default : ch2 = 16'd0;
    endcase

    chan_mix = ch1 + ch2;

    assign sample = chan_mix > 16'hFFFF ? 16'hFFFF : chan_mix[15:0];
  end


endmodule
